module SHA256_tb();

//wire[255:0] t_q; // IHV test
//SHA_IHV dut(.IHV(t_q)); //IHV test
reg t_clk, t_rst;
wire[31:0] t_k;
SHA256_K_machine dut(.clk(t_clk),.rst(t_rst),.K(t_k));
initial 
begin 
//#20 //IHV test
#5
t_clk=0;t_rst=1;
#5
t_clk=1;t_rst=1;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0; t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5
t_clk=1;t_rst=0;
#5
t_clk=0;t_rst=0;
#5


#20
$stop; 
end 

endmodule
